module BCD_7 (
    input wire EN, //��ҳ���ƶ�,EN=0ʱ�ǵ�һҳ��EN=1ʱ�ǵڶ�ҳ
    output reg a,  //���Ϸ���������ܣ���˳ʱ��˳����ת��gΪ�м���������
    output reg b,
    output reg c,
    output reg d,
    output reg e,
    output reg f,
    output reg g
);

    reg [6:0] num;

    always @(*) begin
        if (!EN) begin
            num = 7'b0110000; // ��ʾ����1
        end else begin
            num = 7'b1101101; // ��ʾ����2
        end
        {a, b, c, d, e, f, g} = num;
    end

endmodule
