module control (
    input wire CLK,
    input wire allFull,       // ȫ���ź�
    input wire startWork,     // ��ʼ�������ź�
    output reg isWork         // ����״̬�źţ��ߵ�ƽ��ʾ���ڹ���
);

    always @(posedge CLK) begin
        if (allFull) begin
            // ���ȫ���ź�Ϊ�ߣ�ֹͣ����
            isWork <= 0;
        end else if (startWork) begin
            // �����ʼ�������ź�Ϊ�ߣ���������
            isWork <= 1;
        end
    end

endmodule
